module s();

eqwe

endmodule